module tb_two_bit_adder;

	two_bit_adder tba1(a0, b0, a1, b1, cin0,sum0, sum1, cout1);

	initial begin
	a0 = 0; b0 = 0; a1 = 0; b1 = 0; cin0 = 0; #10;
	a0 = 0; b0 = 0; a1 = 0; b1 = 0; cin0 = 1; #10;
	a0 = 0; b0 = 1; a1 = 0; b1 = 0; cin0 = 0; #10;
	a0 = 1; b0 = 0; a1 = 0; b1 = 0; cin0 = 0; #10;
	a0 = 0; b0 = 1; a1 = 0; b1 = 0; cin0 = 1; #10;
	a0 = 1; b0 = 0; a1 = 0; b1 = 0; cin0 = 1; #10;
	a0 = 1; b0 = 1; a1 = 0; b1 = 0; cin0 = 0; #10;
	a0 = 1; b0 = 1; a1 = 0; b1 = 0; cin0 = 1; #10;
	a0 = 0; b0 = 0; a1 = 0; b1 = 1; cin0 = 0; #10;
	a0 = 0; b0 = 0; a1 = 0; b1 = 1; cin0 = 1; #10;
	a0 = 0; b0 = 1; a1 = 0; b1 = 1; cin0 = 0; #10;
	a0 = 1; b0 = 0; a1 = 0; b1 = 1; cin0 = 0; #10;
	a0 = 0; b0 = 1; a1 = 0; b1 = 1; cin0 = 1; #10;
	a0 = 1; b0 = 0; a1 = 0; b1 = 1; cin0 = 1; #10;
	a0 = 1; b0 = 1; a1 = 0; b1 = 1; cin0 = 0; #10;
	a0 = 1; b0 = 1; a1 = 0; b1 = 1; cin0 = 1; #10;
	a0 = 0; b0 = 0; a1 = 1; b1 = 0; cin0 = 0; #10;
	a0 = 0; b0 = 0; a1 = 1; b1 = 0; cin0 = 1; #10;
	a0 = 0; b0 = 1; a1 = 1; b1 = 0; cin0 = 0; #10;
	a0 = 1; b0 = 0; a1 = 1; b1 = 0; cin0 = 0; #10;
	a0 = 0; b0 = 1; a1 = 1; b1 = 0; cin0 = 1; #10;
	a0 = 1; b0 = 0; a1 = 1; b1 = 0; cin0 = 1; #10;
	a0 = 1; b0 = 1; a1 = 1; b1 = 0; cin0 = 0; #10;
	a0 = 1; b0 = 1; a1 = 1; b1 = 0; cin0 = 1; #10;
	a0 = 0; b0 = 0; a1 = 1; b1 = 1; cin0 = 0; #10;
	a0 = 0; b0 = 0; a1 = 1; b1 = 1; cin0 = 1; #10;
	a0 = 0; b0 = 1; a1 = 1; b1 = 1; cin0 = 0; #10;
	a0 = 1; b0 = 0; a1 = 1; b1 = 1; cin0 = 0; #10;
	a0 = 0; b0 = 1; a1 = 1; b1 = 1; cin0 = 1; #10;
	a0 = 1; b0 = 0; a1 = 1; b1 = 0; cin0 = 1; #10;
	a0 = 1; b0 = 1; a1 = 1; b1 = 1; cin0 = 0; #10;
	a0 = 1; b0 = 1; a1 = 1; b1 = 1; cin0 = 1; #10;
	end
endmodule 