module tb_func;

logic a, b, c, d, f;

func func1 (a, b, c, d, f);


initial begin
	a = 0; b = 0; c = 0; d = 0; #10;
	a = 0; b = 0; c = 0; d = 1; #10;
	a = 0; b = 0; c = 1; d = 0; #10;
	a = 0; b = 0; c = 1; d = 1; #10;
	a = 0; b = 1; c = 0; d = 0; #10;
	a = 0; b = 1; c = 0; d = 1; #10;
	a = 0; b = 1; c = 1; d = 0; #10;
	a = 0; b = 1; c = 1; d = 1; #10;
	a = 1; b = 0; c = 0; d = 0; #10;
	a = 1; b = 0; c = 0; d = 1; #10;
	a = 1; b = 0; c = 1; d = 0; #10;
	a = 1; b = 0; c = 1; d = 1; #10;
	a = 1; b = 1; c = 0; d = 0; #10;
	a = 1; b = 1; c = 0; d = 1; #10;
	a = 1; b = 1; c = 1; d = 0; #10;
	a = 1; b = 1; c = 1; d = 1; #10;
	
end

endmodule	